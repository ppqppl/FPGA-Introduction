module data_drive (input			wire						vga_clk,
                   input			wire						rst_n,
                   input			wire		[ 11:0 ]		addr_h,
                   input			wire		[ 11:0 ]		addr_v,
                   input			wire		[ 2:0 ]		 key,
                   output			reg		[ 15:0 ]				rgb_data);

localparam	red    = 16'd63488;
localparam	orange = 16'd64384;
localparam	yellow = 16'd65472;
localparam	green  = 16'd1024;
localparam	blue   = 16'd31;
localparam	indigo = 16'd18448;
localparam	purple = 16'd32784;
localparam	white  = 16'd65503;
localparam	black  = 16'd0;
reg [ 383:0 ] char_line[ 64:0 ];

localparam	states_1 = 1; // 彩条
localparam	states_2 = 2; // 字符
localparam	states_3 = 3; // 图片

parameter	height = 85; // 图片高度
parameter	width  = 85; // 图片宽度
reg			[ 1:0 ]			states_current			; // 当前状态
reg			[ 1:0 ]			states_next			    ; // 下个状态
reg			[ 13:0 ]		rom_address				; // ROM地址
wire	    [ 15:0 ]		rom_data				; // 图片数据

wire							flag_enable_out1			; // 文字有效区域
wire							flag_enable_out2			; // 图片有效区域
wire							flag_clear_rom_address		; // 地址清零
wire							flag_begin_h			    ; // 图片显示行
wire							flag_begin_v			    ; // 图片显示列

//状态转移
always @( posedge vga_clk or negedge rst_n ) begin
    if ( !rst_n ) begin
        states_current <= states_1;
    end
    else begin
        states_current <= states_next;
    end
end

//状态判断
always @( posedge vga_clk or negedge rst_n ) begin
    if ( !rst_n ) begin
        states_next <= states_1;
    end
    else if ( key[ 0 ] ) begin
        states_next <= states_1;
    end
        else if ( key[ 1 ] ) begin
        states_next <= states_2;
        end
        else if ( key[ 2 ] ) begin
        states_next <= states_3;
        end
    else begin
        states_next <= states_next;
    end
end

//状态输出
always @( * ) begin
    case ( states_current )
        states_1 : begin
            if ( addr_h == 0 ) begin
                rgb_data = black;
            end
            else if ( addr_h >0 && addr_h <81 ) begin
                rgb_data = red;
            end
            else if ( addr_h >80 && addr_h <161 ) begin
                rgb_data = orange;
            end
            else if ( addr_h >160 && addr_h <241 ) begin
                rgb_data = yellow;
            end
            else if ( addr_h >240 && addr_h <321 ) begin
                rgb_data = green;
            end
            else if ( addr_h >320 && addr_h <401 ) begin
                rgb_data = blue;
            end
            else if ( addr_h >400 && addr_h <481 ) begin
                rgb_data = indigo;
            end
            else if ( addr_h >480 && addr_h <561 ) begin
                rgb_data = purple;
            end
            else if ( addr_h >560 && addr_h <641 ) begin
                rgb_data = white;
            end
            else begin
                rgb_data = black;
            end
            
        end
        states_2 : begin
            if ( flag_enable_out1 ) begin
                rgb_data = char_line[ addr_v-208 ][ 532 - addr_h ]? white:black;
            end
            else begin
                rgb_data = black;
            end
        end
        states_3 : begin
            if ( flag_enable_out2 ) begin
                rgb_data = rom_data;
            end
            else begin
                rgb_data = black;
            end
            
        end
        default: begin
            case ( addr_h )
                0 : rgb_data      = black;
                1 : rgb_data      = red;
                81 : rgb_data     = orange;
                161: rgb_data     = yellow;
                241: rgb_data     = green;
                321: rgb_data     = blue;
                401: rgb_data     = indigo;
                481: rgb_data     = purple;
                561: rgb_data     = white;
                default: rgb_data = rgb_data;
            endcase
        end
    endcase
end

assign flag_enable_out1 = states_current == states_2 && addr_h > 148 && addr_h < 533 && addr_v > 208  && addr_v < 273 ;
assign flag_begin_h     = addr_h > ( ( 640 - width ) / 2 ) && addr_h < ( ( 640 - width ) / 2 ) + width + 1;
assign flag_begin_v     = addr_v > ( ( 480 - height )/2 ) && addr_v <( ( 480 - height )/2 ) + height + 1;
assign flag_enable_out2 = states_current == states_3 && flag_begin_h && flag_begin_v;

//ROM地址计数器
always @( posedge vga_clk or negedge rst_n ) begin
    if ( !rst_n ) begin
        rom_address <= 0;
    end
    else if ( flag_clear_rom_address ) begin //计数满清零
        rom_address <= 0;
    end
        else if ( flag_enable_out2 ) begin  //在有效区域内+1
        rom_address <= rom_address + 1;
        end
    else begin  //无效区域保持
        rom_address <= rom_address;
    end
end
assign flag_clear_rom_address = rom_address == height * width - 1;

//初始化显示文字
always@( posedge vga_clk or negedge rst_n ) begin
    if ( !rst_n ) begin
		char_line[0] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[1] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[2] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[3] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[4] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[5] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[6] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[7] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[8] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		char_line[9] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030000000;
		char_line[10] = 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000007F0000000;
		char_line[11] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFF0000000;
		char_line[12] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFF0000000;
		char_line[13] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[14] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[15] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[16] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[17] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[18] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[19] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[20] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[21] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[22] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[23] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[24] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF0000000;
		char_line[25] = 384'h0001C000000000000001C0000000000000000000000000000001C000000000000001C000000000000000000FF0000000;
		char_line[26] = 384'h1FFFC00FFFF000001FFFC00FFFF00000000001FFFC0038001FFFC00FFFF000001FFFC00FFFF000000000000FF0000000;
		char_line[27] = 384'h1FFFC0FFFFFF00001FFFC0FFFFFF000000001FFFFFC0F8001FFFC0FFFFFF00001FFFC0FFFFFF00000000000FF0000000;
		char_line[28] = 384'h003FC3F0003FC000003FC3F0003FC0000000FF0001F1F800003FC3F0003FC000003FC3F0003FC0000000000FF0000000;
		char_line[29] = 384'h001FCF80000FF000001FCF80000FF0000003F800007FF800001FCF80000FF000001FCF80000FF0000000000FF0000000;
		char_line[30] = 384'h001FFE000003FC00001FFE000003FC00000FF000001FF800001FFE000003FC00001FFE000003FC000000000FF0000000;
		char_line[31] = 384'h001FF8000001FE00001FF8000001FE00801FC000000FF800001FF8000001FE00001FF8000001FE000000000FF0000000;
		char_line[32] = 384'h001FE0000000FF00001FE0000000FF00003F80000007F800001FE0000000FF00001FE0000000FF000000000FF0000000;
		char_line[33] = 384'h001FC00000007F00001FC00000007F00007F00000007F800001FC00000007F00001FC00000007F000000000FF0000000;
		char_line[34] = 384'h001FC00000007F80001FC00000007F8000FF00000007F800001FC00000007F80001FC00000007F800000000FF0000000;
		char_line[35] = 384'h001FC00000007F80001FC00000007F8001FE00000007F800001FC00000007F80001FC00000007F800000000FF0000000;
		char_line[36] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[37] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[38] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[39] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[40] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[41] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[42] = 384'h001FC00000003FC0001FC00000003FC001FE00000007F800001FC00000003FC0001FC00000003FC00000000FF0000000;
		char_line[43] = 384'h001FC00000003F80001FC00000003F8001FE00000007F800001FC00000003F80001FC00000003F800000000FF0000000;
		char_line[44] = 384'h001FC00000007F80001FC00000007F8001FE00000007F800001FC00000007F80001FC00000007F800000000FF0000000;
		char_line[45] = 384'h001FC00000007F80001FC00000007F8000FE00000007F800001FC00000007F80001FC00000007F800000000FF0000000;
		char_line[46] = 384'h001FC0000000FF00001FC0000000FF0000FF00000007F800001FC0000000FF00001FC0000000FF000000000FF0000000;
		char_line[47] = 384'h001FC0000001FE00001FC0000001FE00007F00000007F800001FC0000001FE00001FC0000001FE000000000FF0000000;
		char_line[48] = 384'h001FE0000003FC00001FE0000003FC00003F8000000FF800001FE0000003FC00001FE0000003FC000000000FF0000000;
		char_line[49] = 384'h001FF8000007F800001FF8000007F800001FE000001FF800001FF8000007F800001FF8000007F8000000000FF0000000;
		char_line[50] = 384'h001FFC00001FE000001FFC00001FE0000007F000007FF800001FFC00001FE000001FFC00001FE0000000000FF0000000;
		char_line[51] = 384'h001FCF8000FF8000001FCF8000FF80000001FE0007E7F800001FCF8000FF8000001FCF8000FF80000000000FF0000000;
		char_line[52] = 384'h001FC3FFFFFC0000001FC3FFFFFC000000007FFFFF87F800001FC3FFFFFC0000001FC3FFFFFC0000000FFFFFFFFFF000;
		char_line[53] = 384'h001FC03FFFC00000001FC03FFFC00000000007FFF807F800001FC03FFFC00000001FC03FFFC00000000FFFFFFFFFF000;
		char_line[54] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[55] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[56] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[57] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[58] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[59] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[60] = 384'h001FC00000000000001FC00000000000000000000007F800001FC00000000000001FC000000000000000000000000000;
		char_line[61] = 384'h007FF00000000000007FF0000000000000000000000FFE00007FF00000000000007FF000000000000000000000000000;
		char_line[62] = 384'h1FFFFFE0000000001FFFFFE0000000000000000007FFFFF01FFFFFE0000000001FFFFFE0000000000000000000000000;
		char_line[63] = 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
end

//实例化ROM
rom	rom_inst (
.address ( rom_address ),
.clock ( vga_clk ),
.q ( rom_data )
);
endmodule // data_drive

 
 
 
 
 
 
 
 
 
 
 
 
 
