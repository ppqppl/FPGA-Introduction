module uart_driver (
    
);

endmodule //uart_driver