
module Nios (
	clk_clk,
	out_led_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	out_led_export;
	input		reset_reset_n;
endmodule
