// UART.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module UART (
		input  wire       clk_clk,                 //                                clk.clk
		input  wire       reset_reset_n,           //                              reset.reset_n
		input  wire       rs232_0_from_uart_ready, // rs232_0_avalon_data_receive_source.ready
		output wire [7:0] rs232_0_from_uart_data,  //                                   .data
		output wire       rs232_0_from_uart_error, //                                   .error
		output wire       rs232_0_from_uart_valid, //                                   .valid
		input  wire [7:0] rs232_0_to_uart_data,    //  rs232_0_avalon_data_transmit_sink.data
		input  wire       rs232_0_to_uart_error,   //                                   .error
		input  wire       rs232_0_to_uart_valid,   //                                   .valid
		output wire       rs232_0_to_uart_ready,   //                                   .ready
		input  wire       rs232_0_UART_RXD,        //         rs232_0_external_interface.RXD
		output wire       rs232_0_UART_TXD         //                                   .TXD
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> rs232_0:reset

	UART_rs232_0 rs232_0 (
		.clk             (clk_clk),                        //                        clk.clk
		.reset           (rst_controller_reset_out_reset), //                      reset.reset
		.from_uart_ready (rs232_0_from_uart_ready),        // avalon_data_receive_source.ready
		.from_uart_data  (rs232_0_from_uart_data),         //                           .data
		.from_uart_error (rs232_0_from_uart_error),        //                           .error
		.from_uart_valid (rs232_0_from_uart_valid),        //                           .valid
		.to_uart_data    (rs232_0_to_uart_data),           //  avalon_data_transmit_sink.data
		.to_uart_error   (rs232_0_to_uart_error),          //                           .error
		.to_uart_valid   (rs232_0_to_uart_valid),          //                           .valid
		.to_uart_ready   (rs232_0_to_uart_ready),          //                           .ready
		.UART_RXD        (rs232_0_UART_RXD),               //         external_interface.export
		.UART_TXD        (rs232_0_UART_TXD)                //                           .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
