module VGA_String(
OSC_50,     //原CLK2_50时钟信号
VGA_CLK,    //VGA自时钟
VGA_HS,     //行同步信号
VGA_VS,     //场同步信号
VGA_BLANK,  //复合空白信号控制信号  当BLANK为低电平时模拟视频输出消隐电平，此时从R9~R0,G9~G0,B9~B0输入的所有数据被忽略
VGA_SYNC,   //符合同步控制信号      行时序和场时序都要产生同步脉冲
VGA_R,      //VGA绿色
VGA_B,      //VGA蓝色
VGA_G);     //VGA绿色
 input OSC_50;     //外部时钟信号CLK2_50
 output VGA_CLK,VGA_HS,VGA_VS,VGA_BLANK,VGA_SYNC;
 output [7:0] VGA_R,VGA_B,VGA_G;
 parameter H_FRONT = 16;     //行同步前沿信号周期长
 parameter H_SYNC = 96;      //行同步信号周期长
 parameter H_BACK = 48;      //行同步后沿信号周期长
 parameter H_ACT = 640;      //行显示周期长
 parameter H_BLANK = H_FRONT+H_SYNC+H_BACK;        //行空白信号总周期长
 parameter H_TOTAL = H_FRONT+H_SYNC+H_BACK+H_ACT;  //行总周期长耗时
 parameter V_FRONT = 11;     //场同步前沿信号周期长
 parameter V_SYNC = 2;       //场同步信号周期长
 parameter V_BACK = 31;      //场同步后沿信号周期长
 parameter V_ACT = 480;      //场显示周期长
 parameter V_BLANK = V_FRONT+V_SYNC+V_BACK;        //场空白信号总周期长
 parameter V_TOTAL = V_FRONT+V_SYNC+V_BACK+V_ACT;  //场总周期长耗时
 reg [10:0] H_Cont;        //行周期计数器
 reg [10:0] V_Cont;        //场周期计数器
 wire [7:0] VGA_R;         //VGA红色控制线
 wire [7:0] VGA_B;         //VGA绿色控制线
 wire [7:0] VGA_G;         //VGA蓝色控制线
 reg VGA_HS;
 reg VGA_VS;
 reg [10:0] X;             //当前行第几个像素点
 reg [10:0] Y;             //当前场第几行
 reg CLK_25;
 always@(posedge OSC_50)
    begin 
      CLK_25=~CLK_25;         //时钟
    end 
    assign VGA_SYNC = 1'b0;   //同步信号低电平
    assign VGA_BLANK = ~((H_Cont<H_BLANK)||(V_Cont<V_BLANK));  //当行计数器小于行空白总长或场计数器小于场空白总长时，空白信号低电平
    assign VGA_CLK = ~CLK_to_DAC;  //VGA时钟等于CLK_25取反
    assign CLK_to_DAC = CLK_25;
 always@(posedge CLK_to_DAC)
    begin
        if(H_Cont<H_TOTAL)           //如果行计数器小于行总时长
            H_Cont<=H_Cont+1'b1;      //行计数器+1
        else H_Cont<=0;              //否则行计数器清零
        if(H_Cont==H_FRONT-1)        //如果行计数器等于行前沿空白时间-1
            VGA_HS<=1'b0;             //行同步信号置0
        if(H_Cont==H_FRONT+H_SYNC-1) //如果行计数器等于行前沿+行同步-1
            VGA_HS<=1'b1;             //行同步信号置1
        if(H_Cont>=H_BLANK)          //如果行计数器大于等于行空白总时长
            X<=H_Cont-H_BLANK;        //X等于行计数器-行空白总时长   （X为当前行第几个像素点）
        else X<=0;                   //否则X为0
    end
 always@(posedge VGA_HS)
    begin
        if(V_Cont<V_TOTAL)           //如果场计数器小于行总时长
            V_Cont<=V_Cont+1'b1;      //场计数器+1
        else V_Cont<=0;              //否则场计数器清零
        if(V_Cont==V_FRONT-1)       //如果场计数器等于场前沿空白时间-1
            VGA_VS<=1'b0;             //场同步信号置0
        if(V_Cont==V_FRONT+V_SYNC-1) //如果场计数器等于行前沿+场同步-1
            VGA_VS<=1'b1;             //场同步信号置1
        if(V_Cont>=V_BLANK)          //如果场计数器大于等于场空白总时长
            Y<=V_Cont-V_BLANK;        //Y等于场计数器-场空白总时长    （Y为当前场第几行）  
        else Y<=0;                   //否则Y为0
    end
    reg valid_yr;
 always@(posedge CLK_to_DAC)
    if(V_Cont == 10'd56)         //场计数器=32时
        valid_yr<=1'b1;           //行输入激活
    else if(V_Cont==10'd512)     //场计数器=512时
        valid_yr<=1'b0;           //行输入冻结
    wire valid_y=valid_yr;       //连线   
    reg valid_r;            
 always@(posedge CLK_to_DAC)   
    if((H_Cont == 10'd56)&&valid_y)     //行计数器=32时
        valid_r<=1'b1;                   //像素输入激活
    else if((H_Cont==10'd512)&&valid_y) //行计数器=512时 
        valid_r<=1'b0;                   //像素输入冻结
    wire valid = valid_r;               //连线
    wire[10:0] x_dis;     //像素显示控制信号
    wire[10:0] y_dis;     //行显示控制信号
    assign x_dis=X;       //连线X   192 = (640-256 ) /2
    assign y_dis=Y;       //连线Y   231 = (480- 18) /2
        parameter  //点阵字模：每一行char_lineXX是显示的一行，共272列,256
    char_line00=244'h0078000002000000000000000000000000000000000000000000000000000000,  //第1行
    char_line01=244'h27c01ff001000000000000000000000000000000000000000000000000000000,  //第2行
    char_line02=244'h124810107ffe0000000000000000000000000000000000000000000000000000,  //第3行
    char_line03=244'h11501ff04002000018003c003c00180018007e001800180018003c003c003800,  //第4行
    char_line04=244'h87fc101080040000240042004200240024004200240024002400420042004400,  //第5行
    char_line05=244'h41501ff03ff80000400042004200420042000400420040004200420042004200,  //第6行
    char_line06=244'h4248010001000000400002004200420042000400420040004200420042004200,  //第7行
    char_line07=244'h14061100010000005c000400020042004200080042005c004200020002004200,  //第8行
    char_line08=244'h13f81ff801007e00620018000400420042000800420062004200040004004600,  //第9行
    char_line09=244'h22482100fffe0000420004000800420042001000420042004200080008003a00,  //第10行
    char_line0a=244'he248410001000000420002001000420042001000420042004200100010000200,  //第11行
    char_line0b=244'h23f81ff001000000420042002000420042001000420042004200200020000200,  //第12行
    char_line0c=244'h2248010001000000220042004200240024001000240022002400420042002400,  //第13行
    char_line0d=244'h22480100010000001c003c007e0018001800100018001c0018007e007e001800,  //第14行
    char_line0e=244'h23f87ffc05000000000000000000000000000000000000000000000000000000,  //第15行
    char_line0f=244'h0208000002000000000000000000000000000000000000000000000000000000,  //第16行
    char_line10=244'h0000000000000000000000000000000000000000000000000000000000000000,  //第17行
    char_line11=244'h0000000000000000000000000000000000000000000000000000000000000000;  //第18行
    reg [7:0] char_bit;
    always@(posedge CLK_to_DAC)
        if(X==10'd192)char_bit<=8'd256;   //当显示到192像素时准备开始输出图像数据
        else if(X>10'd192&&X<10'd448)     //左边距屏幕192像素到448像素时    448=192+256（图像宽度）
            char_bit<=char_bit-1'b1;       //倒着输出图像信息 
        reg[29:0] VGA_Rgb;                //定义颜色缓存
    always@(posedge CLK_to_DAC)    
        if(X>10'd192&&X<10'd448)    //X控制图像的横向显示边界：左边距屏幕左边192像素  右边界距屏幕左边界448像素
            begin case(Y)            //Y控制图像的纵向显示边界：从距离屏幕顶部200像素开始显示第一行数据
                10'd200:
                if(char_line00[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;  //如果该行有数据 则颜色为红色
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;                      //否则为黑色
                10'd202:
                if(char_line01[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd203:
                if(char_line02[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd204:
                if(char_line03[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd205:
                if(char_line04[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000; 
                10'd206:
                if(char_line05[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd207:
                if(char_line06[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000; 
                10'd208:
                if(char_line07[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd209:
                if(char_line08[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000; 
                10'd210:
                if(char_line09[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd211:
                if(char_line0a[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd212:
                if(char_line0b[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd213:
                if(char_line0c[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd214:
                if(char_line0d[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd215:
                if(char_line0e[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd216:
                if(char_line0f[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd217:
                if(char_line10[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                10'd218:
                if(char_line11[char_bit])VGA_Rgb<=30'b1111111111_0000000000_0000000000;
                else VGA_Rgb<=30'b0000000000_0000000000_0000000000;
                default:VGA_Rgb<=30'h0000000000;   //默认颜色黑色
            endcase 
        end
    else VGA_Rgb<=30'h000000000;             //否则黑色
    assign VGA_R=VGA_Rgb[23:16];
    assign VGA_G=VGA_Rgb[15:8];
    assign VGA_B=VGA_Rgb[7:0];
endmodule



// {010021081110092001003FF8200820083FF8200820083FF82008200820282010},/*"X",0*/

// {04400440044004404444244424481448145014600440044004400440FFFE0000},/*"Y",1*/

// {00007FFC010001001110091009200100FFFE0100010001000100010001000100},/*"P",2*/

// {00000000000000000000000000007FFE00000000000000000000000000000000},/*"-",0*/

// {00000000000007F008181000300037F0380C300C300C300C181807E000000000},/*"6",0*/

// {0000000000000FE0301838180018006001F00018000C380C30180FE000000000},/*"3",1*/

// {00000000000000800780018001800180018001800180018001800FF800000000},/*"1",2*/

// {0000000000000FE03018300C700C301C382C0FCC001C001838300FC000000000},/*"9",3*/

// {00000000000007E01818381C300C300C300C300C300C38181C1007E000000000},/*"0",4*/

// {0000000000001FFC300820100020004000800180030003000380030000000000},/*"7",5*/

// {00000000000007E01818381C300C300C300C300C300C38181C1007E000000000},/*"0",6*/

// {00000000000007F008181000300037F0380C300C300C300C181807E000000000},/*"6",7*/

// {00000000000007E01818381C300C300C300C300C300C38181C1007E000000000},/*"0",8*/

// {0000000000001FF810001000100017F01818000C000C380C30180FE000000000},/*"5",9*/

// {0000000000000FF03018380C101800180060018006000804300C3FF800000000},/*"2",10*/

// {0000000000001FF810001000100017F01818000C000C380C30180FE000000000},/*"5",11*/

