module Nios (
    input  
);
    
endmodule